* NGSPICE file created from cs_flat.ext - technology: sky130A

.subckt cs_flat GND VDS_FR VGS_FR VDD
X0 VDS_FR.t5 VDD.t0 GND sky130_fd_pr__res_xhigh_po_1p41 l=2.12
X1 GND VGS_FR.t0 VDS_FR.t4 GND sky130_fd_pr__nfet_01v8_lvt ad=1.5 pd=6.5 as=1.8 ps=12.6 w=6 l=0.5
X2 GND VGS_FR.t1 VDS_FR.t3 GND sky130_fd_pr__nfet_01v8_lvt ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X3 GND VGS_FR.t2 VDS_FR.t0 GND sky130_fd_pr__nfet_01v8_lvt ad=1.8 pd=12.6 as=1.5 ps=6.5 w=6 l=0.5
X4 VDS_FR.t2 VGS_FR.t3 GND GND sky130_fd_pr__nfet_01v8_lvt ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
X5 VDS_FR.t1 VGS_FR.t4 GND GND sky130_fd_pr__nfet_01v8_lvt ad=1.5 pd=6.5 as=1.5 ps=6.5 w=6 l=0.5
R0 VDS_FR.n5 VDS_FR.n3 256.483
R1 VDS_FR.n21 VDS_FR.n5 185
R2 VDS_FR.n20 VDS_FR.n6 185
R3 VDS_FR.n9 VDS_FR.n7 185
R4 VDS_FR.n16 VDS_FR.n10 185
R5 VDS_FR.n15 VDS_FR.n11 185
R6 VDS_FR.n14 VDS_FR.n12 185
R7 VDS_FR.n13 VDS_FR.t4 180.518
R8 VDS_FR.n6 VDS_FR.n5 144
R9 VDS_FR.n9 VDS_FR.n6 144
R10 VDS_FR.n10 VDS_FR.n9 144
R11 VDS_FR.n11 VDS_FR.n10 144
R12 VDS_FR.n12 VDS_FR.n11 144
R13 VDS_FR.t4 VDS_FR.n12 72.0005
R14 VDS_FR.n22 VDS_FR.n21 27.1064
R15 VDS_FR.n21 VDS_FR.n20 27.1064
R16 VDS_FR.n20 VDS_FR.n7 27.1064
R17 VDS_FR.n16 VDS_FR.n7 27.1064
R18 VDS_FR.n16 VDS_FR.n15 27.1064
R19 VDS_FR.n15 VDS_FR.n14 27.1064
R20 VDS_FR.n24 VDS_FR.n3 25.7837
R21 VDS_FR.n2 VDS_FR.n0 18.4179
R22 VDS_FR.n2 VDS_FR.n1 17.5558
R23 VDS_FR.n23 VDS_FR.n22 9.3005
R24 VDS_FR.n21 VDS_FR.n4 9.3005
R25 VDS_FR.n20 VDS_FR.n19 9.3005
R26 VDS_FR.n18 VDS_FR.n7 9.3005
R27 VDS_FR.n17 VDS_FR.n16 9.3005
R28 VDS_FR.n15 VDS_FR.n8 9.3005
R29 VDS_FR.n22 VDS_FR.n3 9.2683
R30 VDS_FR.n14 VDS_FR.n13 6.30899
R31 VDS_FR.n1 VDS_FR.t3 5.0005
R32 VDS_FR.n1 VDS_FR.t2 5.0005
R33 VDS_FR.n0 VDS_FR.t0 5.0005
R34 VDS_FR.n0 VDS_FR.t1 5.0005
R35 VDS_FR.n25 VDS_FR.n24 4.5005
R36 VDS_FR VDS_FR.t5 3.92989
R37 VDS_FR.n13 VDS_FR.n8 1.21581
R38 VDS_FR.n25 VDS_FR.n2 0.819465
R39 VDS_FR VDS_FR.n25 0.310845
R40 VDS_FR.n23 VDS_FR.n4 0.196152
R41 VDS_FR.n19 VDS_FR.n4 0.196152
R42 VDS_FR.n19 VDS_FR.n18 0.196152
R43 VDS_FR.n18 VDS_FR.n17 0.196152
R44 VDS_FR.n17 VDS_FR.n8 0.196152
R45 VDS_FR.n24 VDS_FR.n23 0.171271
R46 VDD VDD.t0 0.803546
R47 VGS_FR.n2 VGS_FR.t0 486.229
R48 VGS_FR.n0 VGS_FR.t2 486.229
R49 VGS_FR.n2 VGS_FR.t3 485.687
R50 VGS_FR.n1 VGS_FR.t1 485.687
R51 VGS_FR.n0 VGS_FR.t4 485.687
R52 VGS_FR.n1 VGS_FR.n0 0.543978
R53 VGS_FR VGS_FR.n2 0.307565
R54 VGS_FR VGS_FR.n1 0.236913
C0 VDD VDS_FR 0.0934f
C1 VGS_FR VDD 0.00363f
C2 VGS_FR VDS_FR 0.85341f
C3 VGS_FR GND 2.15099f
C4 VDD GND 0.79969f
C5 VDS_FR GND 4.19111f
.ends

