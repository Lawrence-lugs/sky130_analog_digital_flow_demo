* NGSPICE file created from cs_flat.ext - technology: sky130A

.subckt cs_flat GND VDS_FR VDD VGS_FR
X0 GND VGS_FR.t0 VDS_FR.t10 GND sky130_fd_pr__nfet_01v8_lvt ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X1 GND VGS_FR.t1 VDS_FR.t9 GND sky130_fd_pr__nfet_01v8_lvt ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X2 GND VGS_FR.t2 VDS_FR.t8 GND sky130_fd_pr__nfet_01v8_lvt ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X3 VDS_FR.t0 VDD.t0 GND sky130_fd_pr__res_xhigh_po_1p41 l=2.12
X4 GND VGS_FR.t3 VDS_FR.t7 GND sky130_fd_pr__nfet_01v8_lvt ad=0.75 pd=3.5 as=0.9 ps=6.6 w=3 l=0.5
X5 GND VGS_FR.t4 VDS_FR.t6 GND sky130_fd_pr__nfet_01v8_lvt ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X6 VDS_FR.t5 VGS_FR.t5 GND GND sky130_fd_pr__nfet_01v8_lvt ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X7 VDS_FR.t4 VGS_FR.t6 GND GND sky130_fd_pr__nfet_01v8_lvt ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X8 VDS_FR.t3 VGS_FR.t7 GND GND sky130_fd_pr__nfet_01v8_lvt ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X9 VDS_FR.t2 VGS_FR.t8 GND GND sky130_fd_pr__nfet_01v8_lvt ad=0.75 pd=3.5 as=0.75 ps=3.5 w=3 l=0.5
X10 VDS_FR.t1 VGS_FR.t9 GND GND sky130_fd_pr__nfet_01v8_lvt ad=0.9 pd=6.6 as=0.75 ps=3.5 w=3 l=0.5
R0 VGS_FR.n0 VGS_FR.t9 341.63
R1 VGS_FR VGS_FR.t3 341.356
R2 VGS_FR.n7 VGS_FR.t8 341.087
R3 VGS_FR.n6 VGS_FR.t2 341.087
R4 VGS_FR.n5 VGS_FR.t6 341.087
R5 VGS_FR.n4 VGS_FR.t1 341.087
R6 VGS_FR.n3 VGS_FR.t7 341.087
R7 VGS_FR.n2 VGS_FR.t0 341.087
R8 VGS_FR.n1 VGS_FR.t5 341.087
R9 VGS_FR.n0 VGS_FR.t4 341.087
R10 VGS_FR.n1 VGS_FR.n0 0.543978
R11 VGS_FR.n2 VGS_FR.n1 0.543978
R12 VGS_FR.n3 VGS_FR.n2 0.543978
R13 VGS_FR.n4 VGS_FR.n3 0.543978
R14 VGS_FR.n5 VGS_FR.n4 0.543978
R15 VGS_FR.n6 VGS_FR.n5 0.543978
R16 VGS_FR.n7 VGS_FR.n6 0.543978
R17 VGS_FR VGS_FR.n7 0.274957
R18 VDS_FR.n20 VDS_FR.n18 256.483
R19 VDS_FR.n2 VDS_FR.n0 256.483
R20 VDS_FR.n24 VDS_FR.n20 185
R21 VDS_FR.n23 VDS_FR.n21 185
R22 VDS_FR.n6 VDS_FR.n2 185
R23 VDS_FR.n5 VDS_FR.n3 185
R24 VDS_FR.n22 VDS_FR.t7 180.972
R25 VDS_FR.n4 VDS_FR.t1 180.972
R26 VDS_FR.n21 VDS_FR.n20 144
R27 VDS_FR.n3 VDS_FR.n2 144
R28 VDS_FR.t7 VDS_FR.n21 72.0005
R29 VDS_FR.t1 VDS_FR.n3 72.0005
R30 VDS_FR.n17 VDS_FR.n16 29.1983
R31 VDS_FR.n15 VDS_FR.n14 29.1983
R32 VDS_FR.n13 VDS_FR.n12 29.1983
R33 VDS_FR.n11 VDS_FR.n10 29.1983
R34 VDS_FR.n25 VDS_FR.n24 27.1064
R35 VDS_FR.n24 VDS_FR.n23 27.1064
R36 VDS_FR.n7 VDS_FR.n6 27.1064
R37 VDS_FR.n6 VDS_FR.n5 27.1064
R38 VDS_FR.n27 VDS_FR.n18 25.7818
R39 VDS_FR.n9 VDS_FR.n0 25.7818
R40 VDS_FR.n16 VDS_FR.t8 10.0005
R41 VDS_FR.n16 VDS_FR.t2 10.0005
R42 VDS_FR.n14 VDS_FR.t9 10.0005
R43 VDS_FR.n14 VDS_FR.t4 10.0005
R44 VDS_FR.n12 VDS_FR.t10 10.0005
R45 VDS_FR.n12 VDS_FR.t3 10.0005
R46 VDS_FR.n10 VDS_FR.t6 10.0005
R47 VDS_FR.n10 VDS_FR.t5 10.0005
R48 VDS_FR.n26 VDS_FR.n25 9.3005
R49 VDS_FR.n24 VDS_FR.n19 9.3005
R50 VDS_FR.n8 VDS_FR.n7 9.3005
R51 VDS_FR.n6 VDS_FR.n1 9.3005
R52 VDS_FR.n25 VDS_FR.n18 9.2683
R53 VDS_FR.n7 VDS_FR.n0 9.2683
R54 VDS_FR.n23 VDS_FR.n22 6.30296
R55 VDS_FR.n5 VDS_FR.n4 6.30296
R56 VDS_FR.n11 VDS_FR.n9 5.31947
R57 VDS_FR.n28 VDS_FR.n27 4.5005
R58 VDS_FR VDS_FR.t0 3.94993
R59 VDS_FR.n22 VDS_FR.n19 1.22193
R60 VDS_FR.n4 VDS_FR.n1 1.22193
R61 VDS_FR.n13 VDS_FR.n11 0.862569
R62 VDS_FR.n15 VDS_FR.n13 0.862569
R63 VDS_FR.n17 VDS_FR.n15 0.862569
R64 VDS_FR.n28 VDS_FR.n17 0.819465
R65 VDS_FR VDS_FR.n28 0.310845
R66 VDS_FR.n26 VDS_FR.n19 0.196152
R67 VDS_FR.n8 VDS_FR.n1 0.196152
R68 VDS_FR.n27 VDS_FR.n26 0.173988
R69 VDS_FR.n9 VDS_FR.n8 0.173988
R70 VDD VDD.t0 0.803546
C0 VDS_FR VGS_FR 1.10625f
C1 VDD VGS_FR 0.00264f
C2 VDS_FR VDD 0.06853f
C3 VGS_FR GND 3.62596f
C4 VDD GND 0.83505f
C5 VDS_FR GND 5.06078f
.ends

